`timescale 1ns / 1ps
module AL(
    input a;
endmodule
